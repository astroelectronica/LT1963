.title KiCad schematic
.include "C:/AE/LT1963/_models/C3216X5R2A105K160AA_s.mod"
.include "C:/AE/LT1963/_models/CGA5L3X5R1H106K160AB_s.mod"
.include "C:/AE/LT1963/_models/LT1963.lib"
XU3 /VOUT 0 CGA5L3X5R1H106K160AB_s
R2 /VOUT /ADJ {RADJU}
R3 /ADJ 0 {RADJB}
I1 /VOUT 0 {ILOAD}
XU2 /VOUT /ADJ 0 /SHUTDOWN /VIN LT1963
XU1 /VIN 0 C3216X5R2A105K160AA_s
V1 /VIN 0 {VSOURCE}
V2 /SHUTDOWN 0 {VSHDN}
.end
